`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 25.02.2020 11:03:39
// Design Name: 
// Module Name: add_execute
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module add_execute
#(
    parameter len =32
)
(
  input [len-1:0] i_add_pc,
  input [len-1:0] i_shift_sign_extend,
  output [len-1:0] o_add_excute
);

endmodule
