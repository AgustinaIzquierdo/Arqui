`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.11.2019 11:08:40
// Design Name: 
// Module Name: cpu
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`define NB_PC 11
`define NB_OPERANDO 11
`define NB_OPCODE 5
`define RAM_WIDTH 16
`define NB_DECODER_SEL_A 2
`define NB_DECODER 1

module cpu(

    );
endmodule
